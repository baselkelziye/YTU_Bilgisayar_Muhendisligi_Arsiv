module one_bit_xor(out,a,b);
    input a, b;
    output out;

    xor x1(out,a,b);
endmodule


