module one_bit_zeroExtender(out,a);
    input a;
    output out;

    xor(out,a,0);

endmodule


