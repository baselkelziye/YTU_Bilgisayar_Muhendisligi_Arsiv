module one_bit_not(out,a);
    input a;
    output out;

    not n1(out,a);
endmodule


