module one_bit_and(out,a,b);
    input a, b;
    output out;

    and a1(out,a,b);
endmodule


